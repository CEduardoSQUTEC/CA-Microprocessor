module Comparison_part(slt_sel,a,b,result);
    input [31:0] a,b;
    output [31:0] result;
    //Implementar un sign extend

endmodule
