module logic_part()
