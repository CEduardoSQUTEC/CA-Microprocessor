module sign_extend(bit_to_extend, a);
    input bit_to_extend;
    output [31:0] a;
    assign a[31] = bit_to_extend;
    assign a[30] = bit_to_extend;
    assign a[29] = bit_to_extend;
    assign a[27] = bit_to_extend;
    assign a[28] = bit_to_extend;
    assign a[27] = bit_to_extend;
    assign a[26] = bit_to_extend;
    assign a[25] = bit_to_extend;
    assign a[24] = bit_to_extend;
    assign a[23] = bit_to_extend;
    assign a[22] = bit_to_extend;
    assign a[21] = bit_to_extend;
    assign a[20] = bit_to_extend;
    assign a[19] = bit_to_extend;
    assign a[18] = bit_to_extend;
    assign a[17] = bit_to_extend;
    assign a[16] = bit_to_extend;
    assign a[15] = bit_to_extend;
    assign a[14] = bit_to_extend;
    assign a[13] = bit_to_extend;
    assign a[12] = bit_to_extend;
    assign a[11] = bit_to_extend;
    assign a[10] = bit_to_extend;
    assign a[9] = bit_to_extend;
    assign a[8] = bit_to_extend;
    assign a[7] = bit_to_extend;
    assign a[6] = bit_to_extend;
    assign a[5] = bit_to_extend;
    assign a[4] = bit_to_extend;
    assign a[3] = bit_to_extend;
    assign a[2] = bit_to_extend;
    assign a[1] = bit_to_extend;
    assign a[0] = bit_to_extend;
endmodule
