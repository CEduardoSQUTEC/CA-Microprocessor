module arithmetic_part(a,b);
    input a,b;


    
